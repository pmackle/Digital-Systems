module smoothing_filter(

	input [15:0] data_x,
	output [15:0] smooth_out
	
);





endmodule